// baudmux.sv - Baud Divider Mux for UART
// HKL 01 2016

module baudmux
import comm_defs_pkg::*;
(
  input  logic [3:0] baud_sel, // select for baud dividers
  output logic [11:0] baud_div // selected baud divider
);

//---------------------------------------------------------
// Set Baud Rates
//|  SEL | DIV |  10  |  20  |  25  |  30  |  40  |  50  |  60  |  70  |  75  |  80  |  90  | 100  |
//| 4'd0 | 1302|      |      |      |      |      |  9.6K|      |      |      |      |      | 19.2K|
//| 4'd1 |  217|      |      |      |      |      | 57.6K|      |      |      |      |      |115.2K|
//| 4'd2 |  108|      |      | 57.6K|      |      |115.2K|      |      |      |      |      |230.4K|
//| 4'd3 |   54|      |      |115.2K|      |      |230.4K|      |      |      |      |      |460.8K|
//| 4'd4 |   27|      |      |230.4K|      |      |460.8K|      |      |      |      |      |921.6K|
//| 4'd5 |   22|115.2K|230.4K|      |      |460.8K|      |      |      |      |921.6K|      |      |
//| 4'd6 |   20|      |      |      |      |      |      |      |      |921.6K|1.000M|      |      |
//| 4'd7 |   19|      |      |      |      |      |      |      |921.6K|1.000M|      |      |      |
//| 4'd8 |   16|      |      |      |460.8K|      |      |921.6K|      |      |1.250M|      |1.500M|
//| 4'd9 |   15|      |      |      |      |      |      |1.000M|      |1.250M|      |1.500M|      |
//| 4'd10|   10|      |      |      |      |1.000M|1.250M|1.500M|      |      |2.000M|      |      |
//| 4'd11|    8|      |      |      |      |1.250M|1.500M|      |      |      |      |      |3.000M|
//| 4'd12|    6|      |      |1.000M|1.250M|      |2.000M|      |3.000M|3.000M|      |      |      |
//| 4'd13|    5|      |      |1.250M|1.500M|2.000M|      |3.000M|      |      |      |      |      |
//| 4'd14|    4|      |1.250M|1.500M|      |      |3.000M|      |      |      |      |      |      |
//| 4'd15|    2|1.250M|      |3.000M|      |      |      |      |      |      |      |      |      |
//---------------------------------------------------------
always_comb
case(baud_sel)
4'd0 : baud_div = 12'd1302;
4'd1 : baud_div = 12'd217;
4'd2 : baud_div = 12'd108;
4'd3 : baud_div = 12'd54;
4'd4 : baud_div = 12'd27;
4'd5 : baud_div = 12'd22;
4'd6 : baud_div = 12'd20;
4'd7 : baud_div = 12'd19;
4'd8 : baud_div = 12'd16;
4'd9 : baud_div = 12'd15;
4'd10: baud_div = 12'd10;
4'd11: baud_div = 12'd8;
4'd12: baud_div = 12'd6;
4'd13: baud_div = 12'd5;
4'd14: baud_div = 12'd4;
4'd15: baud_div = 12'd2;
default: baud_div = 'x;
endcase

endmodule
